`timescale 1ns / 1ps
module and_gate(i1, i2, d);
	input i1;
	input i2;
	output d;

	// Behaviour design of and2 gate
	// Your code here
	
endmodule
